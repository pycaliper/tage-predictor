../include/common_defines.svh