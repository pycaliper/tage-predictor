`include "common_defines.svh"

module top
    (
        /* verilator lint_off UNUSED */
        input logic clk_i,

        input logic rst_i,

        input logic br_result_i, update_en_i, correct_i,
        input logic [31:0] idx_i,
        /* verilator lint_on UNUSED */
        output logic prediction_o

        , input domain_t domain_i
        , input [31:0] targ_i
        , output logic [31:0] targ_o
    );
    /* verilator lint_off WIDTH */
    //assign prediction_o = `BR_TAKEN;
    //bht b (.*);
    tage_predictor tp (.*);
    /* verilator lint_on WIDTH */
endmodule